library IEEE;
    use IEEE.std_logic_1164.all;
    use IEEE.numeric_std.all;

entity divider is
    port (
        clk: in  std_logic;
        rst: in  std_logic
    );
end entity;

architecture rtl of divider is
begin
end architecture;