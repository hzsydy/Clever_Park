library IEEE;
    use IEEE.std_logic_1164.all;
    use IEEE.numeric_std.all;

entity pwm2int is
    port (
        clk: in  std_logic;
        rst: in  std_logic
    );
end entity;

architecture rtl of pwm2int is
begin
end architecture;